module InstructionMemory(
	input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
);
	always @(*)
		case (Address[11:2])
9'd0: Instruction <= 32'h20100000;
9'd1: Instruction <= 32'h20020014;
9'd2: Instruction <= 32'hac020000;
9'd3: Instruction <= 32'h200241a8;
9'd4: Instruction <= 32'hac020004;
9'd5: Instruction <= 32'h20023af2;
9'd6: Instruction <= 32'hac020008;
9'd7: Instruction <= 32'h3c010000;
9'd8: Instruction <= 32'h3421acda;
9'd9: Instruction <= 32'h00011020;
9'd10: Instruction <= 32'hac02000c;
9'd11: Instruction <= 32'h20020c2b;
9'd12: Instruction <= 32'hac020010;
9'd13: Instruction <= 32'h3c010000;
9'd14: Instruction <= 32'h3421b783;
9'd15: Instruction <= 32'h00011020;
9'd16: Instruction <= 32'hac020014;
9'd17: Instruction <= 32'h3c010000;
9'd18: Instruction <= 32'h3421dac9;
9'd19: Instruction <= 32'h00011020;
9'd20: Instruction <= 32'hac020018;
9'd21: Instruction <= 32'h3c010000;
9'd22: Instruction <= 32'h34218ed9;
9'd23: Instruction <= 32'h00011020;
9'd24: Instruction <= 32'hac02001c;
9'd25: Instruction <= 32'h200209ff;
9'd26: Instruction <= 32'hac020020;
9'd27: Instruction <= 32'h20022f44;
9'd28: Instruction <= 32'hac020024;
9'd29: Instruction <= 32'h2002044e;
9'd30: Instruction <= 32'hac020028;
9'd31: Instruction <= 32'h3c010000;
9'd32: Instruction <= 32'h34219899;
9'd33: Instruction <= 32'h00011020;
9'd34: Instruction <= 32'hac02002c;
9'd35: Instruction <= 32'h20023c56;
9'd36: Instruction <= 32'hac020030;
9'd37: Instruction <= 32'h2002128d;
9'd38: Instruction <= 32'hac020034;
9'd39: Instruction <= 32'h3c010000;
9'd40: Instruction <= 32'h3421dbe3;
9'd41: Instruction <= 32'h00011020;
9'd42: Instruction <= 32'hac020038;
9'd43: Instruction <= 32'h3c010000;
9'd44: Instruction <= 32'h3421d4b4;
9'd45: Instruction <= 32'h00011020;
9'd46: Instruction <= 32'hac02003c;
9'd47: Instruction <= 32'h20023748;
9'd48: Instruction <= 32'hac020040;
9'd49: Instruction <= 32'h20023918;
9'd50: Instruction <= 32'hac020044;
9'd51: Instruction <= 32'h20024112;
9'd52: Instruction <= 32'hac020048;
9'd53: Instruction <= 32'h3c010000;
9'd54: Instruction <= 32'h3421c399;
9'd55: Instruction <= 32'h00011020;
9'd56: Instruction <= 32'hac02004c;
9'd57: Instruction <= 32'h20024955;
9'd58: Instruction <= 32'hac020050;
9'd59: Instruction <= 32'h8c110000;
9'd60: Instruction <= 32'h22270001;
9'd61: Instruction <= 32'h20090004;
9'd62: Instruction <= 32'h222a0000;
9'd63: Instruction <= 32'h20120004;
9'd64: Instruction <= 32'h0c100044;
9'd65: Instruction <= 32'h00000000;
9'd66: Instruction <= 32'hac100000;
9'd67: Instruction <= 32'h08100082;
9'd68: Instruction <= 32'h20080001;
9'd69: Instruction <= 32'h201d0000;
9'd70: Instruction <= 32'hafbf0054;
9'd71: Instruction <= 32'h23bd0004;
9'd72: Instruction <= 32'hac080058;
9'd73: Instruction <= 32'h23bd0004;
9'd74: Instruction <= 32'h0c10005c;
9'd75: Instruction <= 32'h00000000;
9'd76: Instruction <= 32'h23bdfffc;
9'd77: Instruction <= 32'h8c080058;
9'd78: Instruction <= 32'hac08005c;
9'd79: Instruction <= 32'h23bd0004;
9'd80: Instruction <= 32'h0c100070;
9'd81: Instruction <= 32'h00000000;
9'd82: Instruction <= 32'h23bdfffc;
9'd83: Instruction <= 32'h8c08005c;
9'd84: Instruction <= 32'h21080001;
9'd85: Instruction <= 32'h12280002;
9'd86: Instruction <= 32'h08100048;
9'd87: Instruction <= 32'h00000000;
9'd88: Instruction <= 32'h23bdfffc;
9'd89: Instruction <= 32'h8fbf0054;
9'd90: Instruction <= 32'h03e00008;
9'd91: Instruction <= 32'h00000000;
9'd92: Instruction <= 32'h00084880;
9'd93: Instruction <= 32'h01326020;
9'd94: Instruction <= 32'h8d8a0000;
9'd95: Instruction <= 32'h2129fffc;
9'd96: Instruction <= 32'h218cfffc;
9'd97: Instruction <= 32'h22100001;
9'd98: Instruction <= 32'h8d8d0000;
9'd99: Instruction <= 32'h01aa082a;
9'd100: Instruction <= 32'h14200007;
9'd101: Instruction <= 32'h11aa0006;
9'd102: Instruction <= 32'h2129fffc;
9'd103: Instruction <= 32'h218cfffc;
9'd104: Instruction <= 32'h0120082a;
9'd105: Instruction <= 32'h14200002;
9'd106: Instruction <= 32'h08100061;
9'd107: Instruction <= 32'h00000000;
9'd108: Instruction <= 32'h00094882;
9'd109: Instruction <= 32'h212b0001;
9'd110: Instruction <= 32'h03e00008;
9'd111: Instruction <= 32'h00000000;
9'd112: Instruction <= 32'h110b000f;
9'd113: Instruction <= 32'h00084880;
9'd114: Instruction <= 32'h01326020;
9'd115: Instruction <= 32'h000b5080;
9'd116: Instruction <= 32'h8d8b0000;
9'd117: Instruction <= 32'h2129fffc;
9'd118: Instruction <= 32'h218cfffc;
9'd119: Instruction <= 32'h8d8d0000;
9'd120: Instruction <= 32'had8d0004;
9'd121: Instruction <= 32'h2129fffc;
9'd122: Instruction <= 32'h218cfffc;
9'd123: Instruction <= 32'h012a082a;
9'd124: Instruction <= 32'h14200002;
9'd125: Instruction <= 32'h08100077;
9'd126: Instruction <= 32'h00000000;
9'd127: Instruction <= 32'had8b0004;
9'd128: Instruction <= 32'h03e00008;
9'd129: Instruction <= 32'h00000000;
9'd130: Instruction <= 32'h20080000;
9'd131: Instruction <= 32'h1107002e;
9'd132: Instruction <= 32'h200f1d4c;
9'd133: Instruction <= 32'h11e00024;
9'd134: Instruction <= 32'h00084880;
9'd135: Instruction <= 32'h200a0004;
9'd136: Instruction <= 32'h8d2b0000;
9'd137: Instruction <= 32'h1140001d;
9'd138: Instruction <= 32'h200c000f;
9'd139: Instruction <= 32'h018b6024;
9'd140: Instruction <= 32'h20110000;
9'd141: Instruction <= 32'h20120320;
9'd142: Instruction <= 32'h11910004;
9'd143: Instruction <= 32'h22310001;
9'd144: Instruction <= 32'h22520004;
9'd145: Instruction <= 32'h0810008e;
9'd146: Instruction <= 32'h00000000;
9'd147: Instruction <= 32'h8e520000;
9'd148: Instruction <= 32'h200d0004;
9'd149: Instruction <= 32'h01aa6822;
9'd150: Instruction <= 32'h200e0001;
9'd151: Instruction <= 32'h11a00004;
9'd152: Instruction <= 32'h000e7040;
9'd153: Instruction <= 32'h21adffff;
9'd154: Instruction <= 32'h08100097;
9'd155: Instruction <= 32'h00000000;
9'd156: Instruction <= 32'h000e7200;
9'd157: Instruction <= 32'h024e7025;
9'd158: Instruction <= 32'h3c014000;
9'd159: Instruction <= 32'h00200821;
9'd160: Instruction <= 32'hac2e0010;
9'd161: Instruction <= 32'h0c1000ad;
9'd162: Instruction <= 32'h00000000;
9'd163: Instruction <= 32'h000b5902;
9'd164: Instruction <= 32'h214affff;
9'd165: Instruction <= 32'h08100089;
9'd166: Instruction <= 32'h00000000;
9'd167: Instruction <= 32'h21efffff;
9'd168: Instruction <= 32'h08100085;
9'd169: Instruction <= 32'h00000000;
9'd170: Instruction <= 32'h21080001;
9'd171: Instruction <= 32'h08100083;
9'd172: Instruction <= 32'h00000000;
9'd173: Instruction <= 32'h201103e8;
9'd174: Instruction <= 32'h12200003;
9'd175: Instruction <= 32'h2231ffff;
9'd176: Instruction <= 32'h081000ae;
9'd177: Instruction <= 32'h00000000;
9'd178: Instruction <= 32'h03e00008;
9'd179: Instruction <= 32'h00000000;


			default: Instruction <= 32'h00000000;
		endcase
endmodule
